library IEEE; 
use IEEE.STD_LOGIC_1164.all; 


entity DESIGN2TG is 
	port ( 
		BINARY_Y: in STD_LOGIC_VECTOR (8 downto 1); -- 2 Address bits
		MSB_Z: out STD_LOGIC_VECTOR (8 downto 1);
		LSB_Z: out STD_LOGIC_VECTOR (8 downto 1)
	); 
end DESIGN2TG; 

architecture BEHAVIORAL of DESIGN2TG is 
	begin 
	process (BINARY_Y) 

		begin 
		case BINARY_Y is 
			when "01000100" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00000011";--0
			when "01000101" => 
				MSB_Z <="00000011";--0
				LSB_Z <="10011111";--1
			when "01000110" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00100101";--2
			when "01000111" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00001101";--3
			when "01001000" => 
				MSB_Z <="00000011";--0
				LSB_Z <="10011001";--4
			when "01001001" => 
				MSB_Z <="00000011";--0
				LSB_Z <="01001001";--5
			when "01001010" => 
				MSB_Z <="00000011";--0
				LSB_Z <="01000001";--6
			when "01001011" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00011111";--7
			when "01001100" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00000001";--8
			when "01001101" => 
				MSB_Z <="00000011";--0
				LSB_Z <="00001001";--9
			when "01001110" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00000011";--0
			when "01001111" => 
				MSB_Z <="10011111";--1
				LSB_Z <="10011111";--1
			when "01010000" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00100101";--2
			when "01010001" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00001101";--3
			when "01010010" => 
				MSB_Z <="10011111";--1
				LSB_Z <="10011001";--4
			when "01010011" => 
				MSB_Z <="10011111";--1
				LSB_Z <="01001001";--5
			when "01010101" => 
				MSB_Z <="10011111";--1
				LSB_Z <="01000001";--6
			when "01010110" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00011111";--7
			when "01010111" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00000001";--8
			when "01011000" => 
				MSB_Z <="10011111";--1
				LSB_Z <="00001001";--9
			when "01011001" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00000011";--0
			when "01011010" => 
				MSB_Z <="00100101";--2
				LSB_Z <="10011111";--1
			when "01011011" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00100101";--2
			when "01011100" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00001101";--3
			when "01011101" => 
				MSB_Z <="00100101";--2
				LSB_Z <="10011001";--4
			when "01011110" => 
				MSB_Z <="00100101";--2
				LSB_Z <="01001001";--5
			when "01011111" => 
				MSB_Z <="00100101";--2
				LSB_Z <="01000001";--6
			when "01100000" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00011111";--7
			when "01100001" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00000001";--8
			when "01100011" => 
				MSB_Z <="00100101";--2
				LSB_Z <="00001001";--9
			when "01100100" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00000011";--0
			when "01100101" => 
				MSB_Z <="00001101";--3
				LSB_Z <="10011111";--1
			when "01100110" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00100101";--2
			when "01100111" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00001101";--3
			when "01101000" => 
				MSB_Z <="00001101";--3
				LSB_Z <="10011001";--4
			when "01101001" => 
				MSB_Z <="00001101";--3
				LSB_Z <="01001001";--5
			when "01101010" => 
				MSB_Z <="00001101";--3
				LSB_Z <="01000001";--6
			when "01101011" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00011111";--7
			when "01101100" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00000001";--8
			when "01101101" => 
				MSB_Z <="00001101";--3
				LSB_Z <="00001001";--9
			when "01101111" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00000011";--0
			when "01110000" => 
				MSB_Z <="10011001";--4
				LSB_Z <="10011111";--1
			when "01110001" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00100101";--2
			when "01110010" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00001101";--3
			when "01110011" => 
				MSB_Z <="10011001";--4
				LSB_Z <="10011001";--4
			when "01110100" => 
				MSB_Z <="10011001";--4
				LSB_Z <="01001001";--5
			when "01110101" => 
				MSB_Z <="10011001";--4
				LSB_Z <="01000001";--6
			when "01110110" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00011111";--7
			when "01110111" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00000001";--8
			when "01111000" => 
				MSB_Z <="10011001";--4
				LSB_Z <="00001001";--9
			when "01111010" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00000011";--0
			when "01111011" => 
				MSB_Z <="01001001";--5
				LSB_Z <="10011111";--1
			when "01111100" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00100101";--2
			when "01111101" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00001101";--3
			when "01111110" => 
				MSB_Z <="01001001";--5
				LSB_Z <="10011001";--4
			when "01111111" => 
				MSB_Z <="01001001";--5
				LSB_Z <="01001001";--5
			when "10000000" => 
				MSB_Z <="01001001";--5
				LSB_Z <="01000001";--6
			when "10000001" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00011111";--7
			when "10000010" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00000001";--8
			when "10000100" => 
				MSB_Z <="01001001";--5
				LSB_Z <="00001001";--9
			when "10000101" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00000011";--0
			when "10000110" => 
				MSB_Z <="01000001";--6
				LSB_Z <="10011111";--1
			when "10000111" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00100101";--2
			when "10001000" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00001101";--3
			when "10001001" => 
				MSB_Z <="01000001";--6
				LSB_Z <="10011001";--4
			when "10001010" => 
				MSB_Z <="01000001";--6
				LSB_Z <="01001001";--5
			when "10001011" => 
				MSB_Z <="01000001";--6
				LSB_Z <="01000001";--6
			when "10001101" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00011111";--7
			when "10001110" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00000001";--8
			when "10001111" => 
				MSB_Z <="01000001";--6
				LSB_Z <="00001001";--9
			when "10010000" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00000011";--0
			when "10010001" => 
				MSB_Z <="00011111";--7
				LSB_Z <="10011111";--1
			when "10010010" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00100101";--2
			when "10010011" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00001101";--3
			when "10010100" => 
				MSB_Z <="00011111";--7
				LSB_Z <="10011001";--4
			when "10010110" => 
				MSB_Z <="00011111";--7
				LSB_Z <="01001001";--5
			when "10010111" => 
				MSB_Z <="00011111";--7
				LSB_Z <="01000001";--6
			when "10011000" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00011111";--7
			when "10011001" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00000001";--8
			when "10011010" => 
				MSB_Z <="00011111";--7
				LSB_Z <="00001001";--9
			when "10011011" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00000011";--0
			when "10011100" => 
				MSB_Z <="00000001";--8
				LSB_Z <="10011111";--1
			when "10011110" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00100101";--2
			when "10011111" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00001101";--3
			when "10100000" => 
				MSB_Z <="00000001";--8
				LSB_Z <="10011001";--4
			when "10100001" => 
				MSB_Z <="00000001";--8
				LSB_Z <="01001001";--5
			when "10100010" => 
				MSB_Z <="00000001";--8
				LSB_Z <="01000001";--6
			when "10100011" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00011111";--7
			when "10100100" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00000001";--8
			when "10100101" => 
				MSB_Z <="00000001";--8
				LSB_Z <="00001001";--9
			when "10100111" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00000011";--0
			when "10101000" => 
				MSB_Z <="00001001";--9
				LSB_Z <="10011111";--1
			when "10101001" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00100101";--2
			when "10101010" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00001101";--3
			when "10101011" => 
				MSB_Z <="00001001";--9
				LSB_Z <="10011001";--4
			when "10101100" => 
				MSB_Z <="00001001";--9
				LSB_Z <="01001001";--5
			when "10101101" => 
				MSB_Z <="00001001";--9
				LSB_Z <="01000001";--6
			when "10101111" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00011111";--7
			when "10110000" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00000001";--8
			when "10110001" => 
				MSB_Z <="00001001";--9
				LSB_Z <="00001001";--9
			when others => 
				MSB_Z <="10010001";
				LSB_Z <="10010001";
 
		end case; 
	end process; 
end BEHAVIORAL; 
